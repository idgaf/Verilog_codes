module translator(X,H);
	input wire [3:0]X;
	output wire [6:0]H;
	assign H[0]=~X[3]&&~X[2]&&~X[1]&&X[0]||~X[3]&&X[2]&&~X[1]&&~X[0]||X[3]&&~X[2]&&X[1]&&X[0]||X[3]&&X[2]&&~X[1]&&X[0];
	assign H[1]=X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&X[2]&&~X[1]&&X[0]||X[3]&&X[1]&&X[0]||X[2]&&X[1]&&~X[0];
	assign H[2]=X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&~X[2]&&X[1]&&~X[0]||X[3]&&X[2]&&X[1];
	assign H[3]=~X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&~X[2]&&~X[1]&&X[0]||X[2]&&X[1]&&X[0]||X[3]&&~X[2]&&X[1]&&~X[0];
	assign H[4]=~X[3]&&X[2]&&~X[1]||~X[3]&&X[0]||~X[2]&&~X[1]&&X[0];
	assign H[5]=X[3]&&X[2]&&~X[1]&&X[0]||~X[3]&&~X[2]&&X[0]||~X[3]&&X[1]&&X[0]||~X[3]&&~X[2]&&X[1];
	assign H[6]=X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&X[2]&&X[1]&&X[0]||~X[3]&&~X[2]&&~X[1];
endmodule
