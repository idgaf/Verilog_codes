module SuperAdder(a,b,cin,s,cout);
	input wire [3:0]a;
	input wire [3:0]b;
	input wire cin;
	output wire [3:0]s;
	output wire cout;
	wire [3:0]c;
	wire [3:0]G;
	wire [3:0]P;
	assign G[3]=a[3]&&b[3];
	assign G[2]=a[2]&&b[2];
	assign G[1]=a[1]&&b[1];
	assign G[0]=a[0]&&b[0];
	assign P[3]=a[3]&&~b[3]||~a[3]&&b[3];
	assign P[2]=a[2]&&~b[2]||~a[2]&&b[2];
	assign P[1]=a[1]&&~b[1]||~a[1]&&b[1];
	assign P[0]=a[0]&&~b[0]||~a[0]&&b[0];
	wire [3:0]c3;
	wire [2:0]c2;
	wire [1:0]c1;
	and(c3[0],P[3],P[2],P[1],P[0],cin);
	and(c3[1],P[3],P[2],P[1],G[0]);
	and(c3[2],P[3],P[2],G[1]);
	and(c3[3],P[3],G[2]);
	and(c2[0],P[2],P[1],P[0],cin);
	and(c2[1],P[2],P[1],G[0]);
	and(c2[2],P[2],G[1]);
	and(c1[0],P[1],P[0],cin);
	and(c1[1],P[1],G[0]);
	and(c0,P[0],cin);
	or(cout,c3[0],c3[1],c3[2],c3[3],G[3]);
	or(c[2],c2[0],c2[1],c2[2],G[2]);
	or(c[1],c1[0],c1[1],G[1]);
	or(c[0],c0,G[0]);
	assign s[0]=~a[0]&&(~b[0]&&cin||b[0]&&~cin)||a[0]&&(b[0]&&cin||~b[0]&&~cin);
	assign s[1]=~a[1]&&(~b[1]&&c[0]||b[1]&&~c[0])||a[1]&&(b[1]&&c[0]||~b[1]&&~c[0]);
	assign s[2]=~a[2]&&(~b[2]&&c[1]||b[2]&&~c[1])||a[2]&&(b[2]&&c[1]||~b[2]&&~c[1]);
	assign s[3]=~a[3]&&(~b[3]&&c[2]||b[3]&&~c[2])||a[3]&&(b[3]&&c[2]||~b[3]&&~c[2]);
endmodule
	