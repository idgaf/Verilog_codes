`timescale 1ns/1ns
module translator(X,H);
	input [3:0]X;
	output [6:0]H;
	wire [3:0]X;
	wire [6:0]H;
	assign H[0]=~X[3]&&~X[2]&&~X[1]&&X[0]||~X[3]&&X[2]&&~X[1]&&~X[0]||X[3]&&~X[2]&&X[1]&&X[0]||X[3]&&X[2]&&~X[1]&&X[0];
	assign H[1]=X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&X[2]&&~X[1]&&X[0]||X[3]&&X[1]&&X[0]||X[2]&&X[1]&&~X[0];
	assign H[2]=X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&~X[2]&&X[1]&&~X[0]||X[3]&&X[2]&&X[1];
	assign H[3]=~X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&~X[2]&&~X[1]&&X[0]||X[2]&&X[1]&&X[0]||X[3]&&~X[2]&&X[1]&&~X[0];
	assign H[4]=~X[3]&&X[2]&&~X[1]||~X[3]&&X[0]||~X[2]&&~X[1]&&X[0];
	assign H[5]=X[3]&&X[2]&&~X[1]&&X[0]||~X[3]&&~X[2]&&X[0]||~X[3]&&X[1]&&X[0]||~X[3]&&~X[2]&&X[1];
	assign H[6]=X[3]&&X[2]&&~X[1]&&~X[0]||~X[3]&&X[2]&&X[1]&&X[0]||~X[3]&&~X[2]&&~X[1];
endmodule
