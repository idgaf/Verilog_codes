module mux(a,b,s,y);
	input	a,b,s;
	output y;
	wire a,b,s,y;
	assign y=(~s&&a)||(s&&b);
endmodule
