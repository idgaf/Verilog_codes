module Subtractor(A,B,S,sgn);
	input wire [3:0]A;
	input wire [3:0]B;
	output wire [3:0]S;
	output wire sgn;
	wire [3:0]reverse;
	wire [3:0]result;
	wire [3:0]result2;
	assign  reverse = B^(4'b1111);
	wire [3:0]temp;
	RippieAdder (A,reverse,4'b0001,result,sgn);
	assign temp=result^{4{~sgn}};
	RippieAdder (temp,4'b0000,~sgn,S, );
  endmodule