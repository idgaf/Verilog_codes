module postCounter(clk,r,Q);
	input wire clk,r;
	output wire [3:0]Q;
	wire [3:0]self;
	wire [3:0]temp;
	assign self[0]=temp[0];
	assign self[1]=temp[1];
	assign self[2]=temp[2];
	assign self[3]=temp[3];
	DflipflopDescibe a(clk    ,r,temp[0],Q[0],temp[0]);
	DflipflopDescibe b(temp[0],r,temp[1],Q[1],temp[1]);
	DflipflopDescibe c(temp[1],r,temp[2],Q[2],temp[2]);
	DflipflopDescibe d(temp[2],r,temp[3],Q[3],temp[3]);
endmodule

module negCounter(clk,r,Q);
	input wire clk,r;
	output wire [3:0]Q;
	wire [3:0]self;
	wire [3:0]temp;
	assign self[0]=temp[0];
	assign self[1]=temp[1];
	assign self[2]=temp[2];
	assign self[3]=temp[3];
	DflipflopDescibe a(clk ,r,temp[0],Q[0],temp[0]);
	DflipflopDescibe b(Q[0],r,temp[1],Q[1],temp[1]);
	DflipflopDescibe c(Q[1],r,temp[2],Q[2],temp[2]);
	DflipflopDescibe d(Q[2],r,temp[3],Q[3],temp[3]);
endmodule

